package body neorv32_application_image is

constant application_init_image : mem32_t := (
x"000020b7",
x"80008093",
x"30009073",
x"00000097",
x"13808093",
x"30509073",
x"30401073",
x"80000217",
x"3e320213",
x"ff027113",
x"80001197",
x"95c18193",
x"00000293",
x"00000313",
x"00000393",
x"00000413",
x"00000493",
x"00000813",
x"00000893",
x"00000913",
x"00000993",
x"00000a13",
x"00000a93",
x"00000b13",
x"00000b93",
x"00000c13",
x"00000c93",
x"00000d13",
x"00000d93",
x"00000e13",
x"00000e93",
x"00000f13",
x"00000f93",
x"00002597",
x"27c58593",
x"80000617",
x"f7460613",
x"80000697",
x"0f068693",
x"00c58e63",
x"00d65c63",
x"0005a703",
x"00e62023",
x"00458593",
x"00460613",
x"fedff06f",
x"80000717",
x"0cc70713",
x"93818793",
x"00f75863",
x"00072023",
x"00470713",
x"ff5ff06f",
x"00002417",
x"0f040413",
x"00002497",
x"0e848493",
x"00945a63",
x"00042083",
x"000080e7",
x"00440413",
x"ff1ff06f",
x"00000513",
x"00000593",
x"084000ef",
x"30401073",
x"34051073",
x"00000417",
x"03840413",
x"30541073",
x"00002417",
x"0ac40413",
x"00002497",
x"0a448493",
x"00945a63",
x"00042083",
x"000080e7",
x"00440413",
x"ff1ff06f",
x"10500073",
x"ffdff06f",
x"34041073",
x"34202473",
x"01f45413",
x"02041663",
x"34102473",
x"00440413",
x"34141073",
x"34a02473",
x"00347413",
x"ffd40413",
x"00040863",
x"34102473",
x"ffe40413",
x"34141073",
x"34002473",
x"30200073",
x"ff010113",
x"000017b7",
x"00112623",
x"80078793",
x"3047a073",
x"00100593",
x"00100513",
x"7ac000ef",
x"10500073",
x"00000593",
x"00100513",
x"79c000ef",
x"00100593",
x"00300513",
x"790000ef",
x"800e0537",
x"40050513",
x"434000ef",
x"00000593",
x"00300513",
x"778000ef",
x"00100593",
x"00200513",
x"76c000ef",
x"800ca7b7",
x"000366b7",
x"800ca737",
x"af078793",
x"51068693",
x"b1870713",
x"0007a583",
x"00d78633",
x"00478793",
x"00b62023",
x"fee798e3",
x"00000593",
x"00200513",
x"734000ef",
x"00100593",
x"00100513",
x"728000ef",
x"10500073",
x"00000593",
x"00100513",
x"718000ef",
x"00000513",
x"00100593",
x"70c000ef",
x"00c12083",
x"00000513",
x"01010113",
x"00008067",
x"fa010113",
x"02c12023",
x"06412603",
x"06012e83",
x"02e12423",
x"00161713",
x"00f70733",
x"41170733",
x"03d74733",
x"02d12223",
x"40c00633",
x"04812e23",
x"03812e23",
x"04912c23",
x"05212a23",
x"05312823",
x"05412623",
x"05512423",
x"05612223",
x"05712023",
x"03912c23",
x"03a12a23",
x"03b12823",
x"00a12c23",
x"00b12e23",
x"03012623",
x"00060413",
x"00000293",
x"00000f93",
x"03d786b3",
x"00170c13",
x"00d12a23",
x"031886b3",
x"00d12623",
x"02f786b3",
x"02c783b3",
x"00d12823",
x"038fce63",
x"05c12403",
x"05812483",
x"05412903",
x"05012983",
x"04c12a03",
x"04812a83",
x"04412b03",
x"04012b83",
x"03c12c03",
x"03812c83",
x"03412d03",
x"03012d83",
x"06010113",
x"00008067",
x"01812683",
x"00229513",
x"00060593",
x"00a68533",
x"00000493",
x"02412803",
x"00259693",
x"00000a93",
x"00d806b3",
x"00d12423",
x"00000993",
x"00000693",
x"00000b13",
x"00b88d33",
x"02812803",
x"090b5c63",
x"007a8a33",
x"00098913",
x"00000f13",
x"0480006f",
x"00068493",
x"fc1ff06f",
x"01986bb3",
x"000bce63",
x"00fcdc63",
x"00f85a63",
x"000e2b83",
x"00032d83",
x"11bbfbd3",
x"0176f6d3",
x"00180813",
x"004e0e13",
x"00430313",
x"fda81ae3",
x"001f0f13",
x"00fa0a33",
x"01190933",
x"031f5463",
x"00812803",
x"002a1e13",
x"00291313",
x"010e0e33",
x"02c12803",
x"008f0cb3",
x"00680333",
x"00058813",
x"fa1ff06f",
x"00c12803",
x"001b0b13",
x"010989b3",
x"01012803",
x"010a8ab3",
x"f69ff06f",
x"02012803",
x"02080063",
x"01c12803",
x"00082803",
x"0106f6d3",
x"00000813",
x"a1069853",
x"00080463",
x"00000693",
x"00d52023",
x"01d585b3",
x"00148693",
x"00450513",
x"f49714e3",
x"01412683",
x"001f8f93",
x"018282b3",
x"00d383b3",
x"01d40433",
x"ea5ff06f",
x"ffe68793",
x"00200713",
x"02e7c7b3",
x"00000e93",
x"00269693",
x"00000f13",
x"00178793",
x"00279393",
x"00038f93",
x"00fecc63",
x"00008067",
x"00200713",
x"0580006f",
x"00300713",
x"05c0006f",
x"ff010113",
x"00812623",
x"00912423",
x"01212223",
x"00c68433",
x"002f1813",
x"00040893",
x"00062483",
x"00462e03",
x"0008a303",
x"0048a283",
x"a1c49953",
x"00100713",
x"00091663",
x"00048e13",
x"00000713",
x"a06e14d3",
x"fa0496e3",
x"000e0313",
x"a0531e53",
x"fa0e14e3",
x"00030293",
x"d0077753",
x"01050333",
x"00532023",
x"01058333",
x"00e32023",
x"00480813",
x"00860613",
x"00888893",
x"fbf812e3",
x"001e8e93",
x"00ff0f33",
x"007f8fb3",
x"00868633",
x"f8fec2e3",
x"00c12403",
x"00812483",
x"00412903",
x"01010113",
x"00008067",
x"fe010113",
x"01512223",
x"00052a83",
x"00812c23",
x"00912a23",
x"00112e23",
x"01212823",
x"01312623",
x"01412423",
x"00050413",
x"00058493",
x"00100793",
x"0297ce63",
x"00000993",
x"00000a13",
x"0499c863",
x"00000913",
x"06994863",
x"01c12083",
x"01812403",
x"01412483",
x"01012903",
x"00c12983",
x"00812a03",
x"00412a83",
x"02010113",
x"00008067",
x"00279713",
x"00e40733",
x"00072683",
x"a0da96d3",
x"00068463",
x"00072a83",
x"00178793",
x"fa9ff06f",
x"00299913",
x"01240933",
x"00092503",
x"00198993",
x"09557553",
x"3b8000ef",
x"00a92023",
x"00092783",
x"00fa7a53",
x"f8dff06f",
x"00291993",
x"013409b3",
x"0009a503",
x"000a0593",
x"00190913",
x"4e1000ef",
x"00a9a023",
x"f75ff06f",
x"fc010113",
x"02812c23",
x"02912a23",
x"03212823",
x"03412423",
x"80000437",
x"ffff6a37",
x"7ff89937",
x"800004b7",
x"03312623",
x"03512223",
x"03612023",
x"01712e23",
x"01812c23",
x"02112e23",
x"00050993",
x"65840413",
x"01900c13",
x"568a0a13",
x"31000b93",
x"68090913",
x"00200b13",
x"00100a93",
x"67048493",
x"03840833",
x"00040593",
x"01612223",
x"01512023",
x"00500893",
x"01c00793",
x"00100713",
x"00098693",
x"00100613",
x"03740533",
x"01480833",
x"00440413",
x"01250533",
x"bc5ff0ef",
x"fc9414e3",
x"800c5437",
x"7fdad9b7",
x"00001937",
x"800c64b7",
x"d8040413",
x"e0098993",
x"26090913",
x"fe048493",
x"00241613",
x"012405b3",
x"00040513",
x"01c00693",
x"01360633",
x"31040413",
x"d79ff0ef",
x"fe9412e3",
x"80003437",
x"7fe64a37",
x"7ffb5937",
x"800c59b7",
x"800034b7",
x"bf040413",
x"09600b93",
x"7d0a0a13",
x"06400b13",
x"88090913",
x"00100a93",
x"d8098993",
x"c3048493",
x"03740833",
x"00040593",
x"00012223",
x"01512023",
x"00500893",
x"00e00793",
x"00600713",
x"00098693",
x"00100613",
x"03640533",
x"01480833",
x"00440413",
x"01250533",
x"b15ff0ef",
x"fc9414e3",
x"800c9437",
x"7fda4937",
x"800c94b7",
x"b4040413",
x"54090913",
x"18048493",
x"00241613",
x"64040593",
x"00040513",
x"00a00693",
x"01260633",
x"06440413",
x"cd1ff0ef",
x"fe9412e3",
x"800c97b7",
x"ec468537",
x"800c9837",
x"fff688b7",
x"800ca637",
x"7c078793",
x"00000593",
x"19000e13",
x"4f050513",
x"18080813",
x"27088893",
x"9a060613",
x"03c78333",
x"800c9737",
x"00b7a023",
x"b4070713",
x"00a30333",
x"00e306b3",
x"0006a683",
x"00072f03",
x"0007ae83",
x"00470713",
x"11e6f6d3",
x"01d6f6d3",
x"00d7a023",
x"ff0710e3",
x"01178733",
x"00072683",
x"0007a703",
x"00d77753",
x"00e7a023",
x"0007a703",
x"a0b71753",
x"00070463",
x"00b7a023",
x"00478793",
x"fac790e3",
x"fa0e8537",
x"800ca837",
x"fff728b7",
x"800ca637",
x"00000593",
x"07800e13",
x"15050513",
x"9a080813",
x"ff088893",
x"af060613",
x"03c78333",
x"800c9737",
x"00b7a023",
x"7c070713",
x"00a30333",
x"00e306b3",
x"0006a683",
x"00072f03",
x"0007ae83",
x"00470713",
x"11e6f6d3",
x"01d6f6d3",
x"00d7a023",
x"ff0710e3",
x"011786b3",
x"0006a303",
x"0007a683",
x"0066f6d3",
x"00d7a023",
x"0007a683",
x"a0b696d3",
x"00068463",
x"00b7a023",
x"00478793",
x"fac790e3",
x"fbd45837",
x"800ca8b7",
x"fff735b7",
x"800ca637",
x"00000e13",
x"05400e93",
x"a8080813",
x"af088893",
x"d1058593",
x"b1860613",
x"03d78333",
x"01c7a023",
x"00070513",
x"01030333",
x"00a306b3",
x"0006a683",
x"00052f83",
x"0007af03",
x"00450513",
x"11f6f6d3",
x"01e6f6d3",
x"00d7a023",
x"ff1510e3",
x"00b786b3",
x"0006a303",
x"0007a683",
x"00478793",
x"0066f6d3",
x"fed7ae23",
x"fac79ae3",
x"03812403",
x"03c12083",
x"03412483",
x"03012903",
x"02c12983",
x"02812a03",
x"02412a83",
x"02012b03",
x"01c12b83",
x"01812c03",
x"00a00593",
x"04010113",
x"be1ff06f",
x"00100793",
x"00a797b3",
x"02052513",
x"00154513",
x"00251513",
x"c0852703",
x"00058863",
x"00f767b3",
x"c0f52423",
x"00008067",
x"fff7c793",
x"00e7f7b3",
x"ff1ff06f",
x"ff010113",
x"00812423",
x"00912223",
x"00112623",
x"00050413",
x"0a8000ef",
x"00050493",
x"00040513",
x"088000ef",
x"02050663",
x"800007b7",
x"1247a583",
x"00040513",
x"4a1000ef",
x"02a04863",
x"800007b7",
x"1287a583",
x"00040513",
x"539000ef",
x"04054463",
x"00c12083",
x"00812403",
x"00048513",
x"00412483",
x"01010113",
x"00008067",
x"4bc000ef",
x"800007b7",
x"1207a483",
x"00c12083",
x"00812403",
x"02200793",
x"00f52023",
x"00048513",
x"00412483",
x"01010113",
x"00008067",
x"490000ef",
x"02200793",
x"00f52023",
x"00000493",
x"fadff06f",
x"00151513",
x"7f8007b7",
x"00155513",
x"00f52533",
x"00008067",
x"fe010113",
x"00151793",
x"00812c23",
x"00112e23",
x"0017d793",
x"7f800737",
x"00050413",
x"18f76863",
x"01212823",
x"01f55913",
x"2ae78e63",
x"42b17737",
x"21770713",
x"26a74a63",
x"28054463",
x"3eb17737",
x"00912a23",
x"01312623",
x"21870713",
x"16f77c63",
x"3f851737",
x"01412423",
x"01512223",
x"59170713",
x"2ef76a63",
x"800007b7",
x"00291493",
x"17078793",
x"009787b3",
x"0007a583",
x"00040513",
x"040010ef",
x"800007b7",
x"16878793",
x"009787b3",
x"0007aa83",
x"00194493",
x"00050993",
x"412484b3",
x"000a8593",
x"00098513",
x"018010ef",
x"00050593",
x"00050413",
x"4c1000ef",
x"800007b7",
x"1387a583",
x"00050913",
x"4b1000ef",
x"800007b7",
x"13c7a583",
x"7f1000ef",
x"00090593",
x"49d000ef",
x"800007b7",
x"1407a583",
x"394000ef",
x"00090593",
x"489000ef",
x"800007b7",
x"1447a583",
x"7c9000ef",
x"00090593",
x"475000ef",
x"800007b7",
x"1487a583",
x"36c000ef",
x"00090593",
x"461000ef",
x"00050593",
x"00040513",
x"7a1000ef",
x"00050593",
x"00050913",
x"00040513",
x"445000ef",
x"00050a13",
x"28048a63",
x"800007b7",
x"1547a503",
x"00090593",
x"779000ef",
x"00050593",
x"000a0513",
x"744000ef",
x"00050593",
x"000a8513",
x"761000ef",
x"00098593",
x"759000ef",
x"800007b7",
x"00050593",
x"1507a503",
x"749000ef",
x"f8300793",
x"16f4ce63",
x"01749493",
x"00a48533",
x"01c12083",
x"01812403",
x"01412483",
x"01012903",
x"00c12983",
x"00812a03",
x"00412a83",
x"02010113",
x"00008067",
x"00050593",
x"2c4000ef",
x"01c12083",
x"01812403",
x"02010113",
x"00008067",
x"34000737",
x"14e7e663",
x"800009b7",
x"00040593",
x"00040513",
x"399000ef",
x"800007b7",
x"1387a583",
x"00050493",
x"389000ef",
x"800007b7",
x"13c7a583",
x"6c9000ef",
x"00048593",
x"375000ef",
x"800007b7",
x"1407a583",
x"26c000ef",
x"00048593",
x"361000ef",
x"800007b7",
x"1447a583",
x"6a1000ef",
x"00048593",
x"34d000ef",
x"800007b7",
x"1487a583",
x"244000ef",
x"00048593",
x"339000ef",
x"00050593",
x"00040513",
x"679000ef",
x"00050913",
x"00090593",
x"00040513",
x"31d000ef",
x"800007b7",
x"1547a583",
x"00050493",
x"00090513",
x"655000ef",
x"00050593",
x"00048513",
x"620000ef",
x"00040593",
x"641000ef",
x"00050593",
x"1509a503",
x"635000ef",
x"01c12083",
x"01812403",
x"01412483",
x"01012903",
x"00c12983",
x"02010113",
x"00008067",
x"01812403",
x"01012903",
x"01c12083",
x"00000513",
x"02010113",
x"1a00006f",
x"42cff737",
x"1b570713",
x"d6f77ae3",
x"01812403",
x"01012903",
x"01c12083",
x"00000513",
x"02010113",
x"1700006f",
x"00000513",
x"0c091c63",
x"01012903",
x"00040513",
x"ec1ff06f",
x"800007b7",
x"1587a583",
x"06448493",
x"01749493",
x"00a48533",
x"265000ef",
x"e79ff06f",
x"800007b7",
x"14c7a583",
x"00040513",
x"800009b7",
x"150000ef",
x"1509a483",
x"00048593",
x"0e9000ef",
x"e8a05ee3",
x"00048593",
x"00040513",
x"134000ef",
x"01412483",
x"01012903",
x"00c12983",
x"e65ff06f",
x"800007b7",
x"12c7a583",
x"00040513",
x"00291913",
x"20d000ef",
x"800007b7",
x"17878793",
x"012787b3",
x"0007a583",
x"0fc000ef",
x"170010ef",
x"00050493",
x"1d8010ef",
x"800007b7",
x"1307a583",
x"00050913",
x"1dd000ef",
x"00050593",
x"00040513",
x"51d000ef",
x"800007b7",
x"1347a583",
x"00050993",
x"00090513",
x"1bd000ef",
x"00050a93",
x"ce1ff06f",
x"01012903",
x"df1ff06f",
x"00812a03",
x"00412a83",
x"800009b7",
x"e79ff06f",
x"ff010113",
x"00812423",
x"00912223",
x"00112623",
x"00050413",
x"00058493",
x"078000ef",
x"00952023",
x"00c12083",
x"00040513",
x"00812403",
x"00412483",
x"01010113",
x"00008067",
x"ff010113",
x"00112623",
x"02050063",
x"80000537",
x"00b54533",
x"14d000ef",
x"00c12083",
x"02200593",
x"01010113",
x"fa5ff06f",
x"00058513",
x"135000ef",
x"00c12083",
x"02200593",
x"01010113",
x"f8dff06f",
x"800007b7",
x"15c7a583",
x"fb9ff06f",
x"800007b7",
x"1607a583",
x"fadff06f",
x"800007b7",
x"1807a503",
x"00008067",
x"008006b7",
x"fff68693",
x"ff010113",
x"00a6f633",
x"01755713",
x"00812423",
x"01f55413",
x"00361513",
x"0175d613",
x"00b6f6b3",
x"01212023",
x"0ff67613",
x"0ff77913",
x"00112623",
x"00912223",
x"01f5d593",
x"00369793",
x"40c906b3",
x"18b41063",
x"08d05c63",
x"02061663",
x"02078063",
x"fff90693",
x"00069863",
x"00a787b3",
x"00100913",
x"04c0006f",
x"0ff00713",
x"00e91e63",
x"00050793",
x"10c0006f",
x"0ff00713",
x"fee90ae3",
x"04000737",
x"00e7e7b3",
x"01b00613",
x"00100713",
x"00d64e63",
x"02000613",
x"00d7d733",
x"40d606b3",
x"00d796b3",
x"00d036b3",
x"00d76733",
x"00a707b3",
x"00579713",
x"0c075663",
x"00190913",
x"0ff00713",
x"2ce90a63",
x"7e000737",
x"0017f693",
x"fff70713",
x"0017d793",
x"00e7f7b3",
x"00d7e7b3",
x"0a40006f",
x"06068663",
x"41260733",
x"02091063",
x"0c050863",
x"fff70693",
x"f60684e3",
x"0ff00593",
x"02b71063",
x"0ff00913",
x"07c0006f",
x"0ff00693",
x"fed60ae3",
x"040006b7",
x"00d56533",
x"00070693",
x"01b00593",
x"00100713",
x"00d5ce63",
x"02000713",
x"40d70733",
x"00e51733",
x"00d555b3",
x"00e03733",
x"00e5e733",
x"00e787b3",
x"00060913",
x"f69ff06f",
x"00190713",
x"0fe77693",
x"04069c63",
x"04091263",
x"02050263",
x"f00788e3",
x"00a787b3",
x"00579713",
x"00075a63",
x"fc000737",
x"fff70713",
x"00e7f7b3",
x"00100913",
x"0077f713",
x"20070a63",
x"00f7f713",
x"00400693",
x"20d70463",
x"00478793",
x"2000006f",
x"f60502e3",
x"16079663",
x"00050793",
x"f59ff06f",
x"0ff00693",
x"1ed70063",
x"00f507b3",
x"0017d793",
x"00070913",
x"fc1ff06f",
x"06d05e63",
x"06061263",
x"ea0782e3",
x"fff90693",
x"00069863",
x"40f507b3",
x"00100913",
x"0340006f",
x"0ff00713",
x"e8e904e3",
x"01b00613",
x"00100713",
x"00d64e63",
x"02000613",
x"00d7d733",
x"40d606b3",
x"00d796b3",
x"00d036b3",
x"00d76733",
x"40e507b3",
x"00579713",
x"f60754e3",
x"040004b7",
x"fff48493",
x"0097f4b3",
x"1080006f",
x"0ff00713",
x"e4e900e3",
x"04000737",
x"00e7e7b3",
x"fb1ff06f",
x"06068e63",
x"41260733",
x"02091663",
x"1a050e63",
x"fff70693",
x"00069863",
x"40a787b3",
x"00058413",
x"f7dff06f",
x"0ff00813",
x"03071063",
x"0ff00913",
x"19c0006f",
x"0ff00693",
x"fed60ae3",
x"040006b7",
x"00d56533",
x"00070693",
x"01b00813",
x"00100713",
x"00d84e63",
x"02000713",
x"40d70733",
x"00e51733",
x"00d55833",
x"00e03733",
x"00e86733",
x"40e787b3",
x"00060913",
x"00058413",
x"f5dff06f",
x"00190713",
x"0fe77713",
x"04071c63",
x"02091c63",
x"00051863",
x"12079e63",
x"00000413",
x"0c00006f",
x"d8078ae3",
x"40f50733",
x"00571693",
x"40a787b3",
x"1206c063",
x"00070793",
x"e80716e3",
x"00000793",
x"fd9ff06f",
x"ea0510e3",
x"00058413",
x"de079ce3",
x"00000413",
x"020007b7",
x"0ff00913",
x"0800006f",
x"40f504b3",
x"00549713",
x"04075463",
x"40a784b3",
x"00058413",
x"00048513",
x"791000ef",
x"ffb50513",
x"00a494b3",
x"03254e63",
x"41250533",
x"00150513",
x"02000713",
x"40a70733",
x"00a4d7b3",
x"00e494b3",
x"009034b3",
x"0097e7b3",
x"00000913",
x"e19ff06f",
x"fc0492e3",
x"00000793",
x"00000913",
x"f5dff06f",
x"fc0007b7",
x"fff78793",
x"40a90933",
x"00f4f7b3",
x"df5ff06f",
x"0ff00913",
x"00000793",
x"00579713",
x"00075e63",
x"00190913",
x"0ff00713",
x"06e90663",
x"fc000737",
x"fff70713",
x"00e7f7b3",
x"0ff00713",
x"0037d793",
x"00e91863",
x"00078663",
x"004007b7",
x"00000413",
x"00c12083",
x"01791713",
x"01f41513",
x"7f8006b7",
x"00812403",
x"00979793",
x"00d77733",
x"0097d793",
x"00f767b3",
x"00412483",
x"00012903",
x"00a7e533",
x"01010113",
x"00008067",
x"00070913",
x"00058413",
x"d71ff06f",
x"00000793",
x"fa1ff06f",
x"fd010113",
x"02912223",
x"01755493",
x"01312e23",
x"01512a23",
x"01612823",
x"00951a93",
x"02112623",
x"02812423",
x"03212023",
x"01412c23",
x"01712623",
x"01812423",
x"0ff4f493",
x"00058b13",
x"009ada93",
x"01f55993",
x"08048463",
x"0ff00793",
x"0af48063",
x"003a9a93",
x"040007b7",
x"00faeab3",
x"f8148493",
x"00000b93",
x"017b5793",
x"009b1413",
x"0ff7f793",
x"00945413",
x"01fb5b13",
x"08078a63",
x"0ff00713",
x"0ae78663",
x"00341413",
x"04000737",
x"00e46433",
x"f8178793",
x"00000713",
x"40f48a33",
x"002b9793",
x"00e7e7b3",
x"fff78793",
x"00e00693",
x"0169c933",
x"08f6ee63",
x"000026b7",
x"00279793",
x"1c468693",
x"00d787b3",
x"0007a783",
x"00078067",
x"020a8a63",
x"000a8513",
x"5d5000ef",
x"ffb50793",
x"f8a00493",
x"00fa9ab3",
x"40a484b3",
x"f79ff06f",
x"0ff00493",
x"00200b93",
x"f60a88e3",
x"00300b93",
x"f69ff06f",
x"00000493",
x"00100b93",
x"f5dff06f",
x"02040a63",
x"00040513",
x"595000ef",
x"ffb50793",
x"00f41433",
x"f8a00793",
x"40a787b3",
x"f6dff06f",
x"0ff00793",
x"00200713",
x"f60402e3",
x"00300713",
x"f5dff06f",
x"00000793",
x"00100713",
x"f51ff06f",
x"00541c13",
x"168af863",
x"fffa0a13",
x"00000413",
x"010c5b13",
x"000109b7",
x"000b0593",
x"fe098993",
x"000a8513",
x"48d000ef",
x"013c79b3",
x"00050593",
x"00050b93",
x"00098513",
x"44d000ef",
x"00050493",
x"000b0593",
x"000a8513",
x"4b1000ef",
x"01045793",
x"01051513",
x"00a7e7b3",
x"000b8413",
x"0097fe63",
x"00fc07b3",
x"fffb8413",
x"0187e863",
x"0097f663",
x"ffeb8413",
x"018787b3",
x"409784b3",
x"000b0593",
x"00048513",
x"42d000ef",
x"00050593",
x"00050a93",
x"00098513",
x"3f1000ef",
x"00050993",
x"000b0593",
x"00048513",
x"455000ef",
x"01051793",
x"000a8713",
x"0337f263",
x"018786b3",
x"00f6b633",
x"fffa8713",
x"00068793",
x"00061863",
x"0136f663",
x"ffea8713",
x"018687b3",
x"01041413",
x"413787b3",
x"00e46433",
x"00f037b3",
x"00f46433",
x"07fa0713",
x"0ce05e63",
x"00747793",
x"00078a63",
x"00f47793",
x"00400693",
x"00d78463",
x"00440413",
x"00441793",
x"0007da63",
x"f80007b7",
x"fff78793",
x"00f47433",
x"080a0713",
x"0fe00793",
x"08e7c063",
x"00345793",
x"02c12083",
x"02812403",
x"00979793",
x"01771713",
x"0097d793",
x"01f91513",
x"00f76733",
x"02412483",
x"02012903",
x"01c12983",
x"01812a03",
x"01412a83",
x"01012b03",
x"00c12b83",
x"00812c03",
x"00a76533",
x"03010113",
x"00008067",
x"01fa9413",
x"001ada93",
x"e95ff06f",
x"00098913",
x"000a8413",
x"000b8713",
x"00300793",
x"08f70663",
x"00100793",
x"08f70a63",
x"00200793",
x"f4f714e3",
x"00000793",
x"0ff00713",
x"f81ff06f",
x"000b0913",
x"fd9ff06f",
x"00400437",
x"00000913",
x"00300713",
x"fc9ff06f",
x"00100793",
x"40e787b3",
x"01b00713",
x"04f74c63",
x"09ea0493",
x"00f457b3",
x"00941433",
x"00803433",
x"0087e7b3",
x"0077f713",
x"00070a63",
x"00f7f713",
x"00400693",
x"00d70463",
x"00478793",
x"00579713",
x"0037d793",
x"02075263",
x"00000793",
x"00100713",
x"f15ff06f",
x"004007b7",
x"0ff00713",
x"00000913",
x"f05ff06f",
x"00000793",
x"00000713",
x"ef9ff06f",
x"008007b7",
x"fff78793",
x"01755693",
x"00a7f633",
x"01f55713",
x"0ff6f693",
x"0175d513",
x"0ff00813",
x"00b7f7b3",
x"0ff57513",
x"01f5d593",
x"01069463",
x"04061263",
x"0ff00813",
x"01051463",
x"02079c63",
x"04069a63",
x"02051c63",
x"04061863",
x"04078263",
x"00100513",
x"02059e63",
x"fff00513",
x"00008067",
x"fea6c8e3",
x"02c7e263",
x"00000513",
x"02f67263",
x"fe1ff06f",
x"ffe00513",
x"00008067",
x"fc060ae3",
x"00e59e63",
x"fcd55ee3",
x"fff00513",
x"00058c63",
x"00008067",
x"fe0516e3",
x"fe0794e3",
x"fff00513",
x"fe0718e3",
x"00100513",
x"00008067",
x"008007b7",
x"fff78793",
x"01755693",
x"00a7f633",
x"01f55713",
x"0ff6f693",
x"0175d513",
x"0ff00813",
x"00b7f7b3",
x"0ff57513",
x"01f5d593",
x"01069463",
x"04061263",
x"0ff00813",
x"01051463",
x"02079c63",
x"04069a63",
x"02051c63",
x"04061863",
x"04078263",
x"00100513",
x"02059e63",
x"fff00513",
x"00008067",
x"fea6c8e3",
x"02c7e263",
x"00000513",
x"02f67263",
x"fe1ff06f",
x"00200513",
x"00008067",
x"fc060ae3",
x"00e59e63",
x"fcd55ee3",
x"fff00513",
x"00058c63",
x"00008067",
x"fe0516e3",
x"fe0794e3",
x"fff00513",
x"fe0718e3",
x"00100513",
x"00008067",
x"fe010113",
x"01212823",
x"01755913",
x"00912a23",
x"01312623",
x"01512223",
x"00951493",
x"00112e23",
x"00812c23",
x"01412423",
x"0ff97913",
x"00058a93",
x"0094d493",
x"01f55993",
x"14090063",
x"0ff00793",
x"14f90c63",
x"00349493",
x"040007b7",
x"00f4e4b3",
x"f8190913",
x"00000a13",
x"017ad793",
x"009a9413",
x"0ff7f793",
x"00945413",
x"01fada93",
x"14078663",
x"0ff00713",
x"16e78263",
x"00341413",
x"04000737",
x"00e46433",
x"f8178793",
x"00000713",
x"00f90933",
x"002a1793",
x"00e7e7b3",
x"00a00693",
x"00190813",
x"20f6ca63",
x"00200693",
x"0159c9b3",
x"14f6c663",
x"fff78793",
x"00100693",
x"16f6f263",
x"00010eb7",
x"fffe8313",
x"0104df13",
x"01045793",
x"0064f4b3",
x"00647433",
x"00048513",
x"00040593",
x"019000ef",
x"00050893",
x"00078593",
x"00048513",
x"009000ef",
x"00050713",
x"00040593",
x"000f0513",
x"7f8000ef",
x"00050e13",
x"00078593",
x"000f0513",
x"7e8000ef",
x"0108d793",
x"01c70733",
x"00e787b3",
x"00050693",
x"01c7f463",
x"01d506b3",
x"0067f733",
x"01071713",
x"0068f8b3",
x"01170733",
x"0107d793",
x"00671413",
x"00d787b3",
x"01a75713",
x"00679793",
x"00803433",
x"00e46433",
x"00479713",
x"0087e433",
x"00075a63",
x"00145793",
x"00147413",
x"0087e433",
x"00080913",
x"00090813",
x"0c00006f",
x"02048a63",
x"00048513",
x"04d000ef",
x"ffb50793",
x"f8a00913",
x"00f494b3",
x"40a90933",
x"ec1ff06f",
x"0ff00913",
x"00200a13",
x"ea048ce3",
x"00300a13",
x"eb1ff06f",
x"00000913",
x"00100a13",
x"ea5ff06f",
x"02040a63",
x"00040513",
x"00d000ef",
x"ffb50793",
x"00f41433",
x"f8a00793",
x"40a787b3",
x"eb5ff06f",
x"0ff00793",
x"00200713",
x"ea0406e3",
x"00300713",
x"ea5ff06f",
x"00000793",
x"00100713",
x"e99ff06f",
x"00100693",
x"00f697b3",
x"5307f693",
x"0c069063",
x"2407f693",
x"12069263",
x"0887f793",
x"ea0784e3",
x"000a8993",
x"00200793",
x"10f70263",
x"00300793",
x"10f70463",
x"00100793",
x"10f70863",
x"07f80713",
x"08e05c63",
x"00747793",
x"00078a63",
x"00f47793",
x"00400693",
x"00d78463",
x"00440413",
x"00441793",
x"0007da63",
x"f80007b7",
x"fff78793",
x"00f47433",
x"08080713",
x"0fe00793",
x"0ae7ca63",
x"00345793",
x"01c12083",
x"01812403",
x"00979793",
x"01771513",
x"0097d793",
x"01f99993",
x"00f56533",
x"01412483",
x"01012903",
x"00812a03",
x"00412a83",
x"01356533",
x"00c12983",
x"02010113",
x"00008067",
x"00f00693",
x"06d78c63",
x"00b00693",
x"f4d78ce3",
x"00048413",
x"000a0713",
x"f51ff06f",
x"00100793",
x"40e787b3",
x"01b00713",
x"06f74263",
x"09e80813",
x"01041833",
x"00f457b3",
x"01003833",
x"0107e7b3",
x"0077f713",
x"00070a63",
x"00f7f713",
x"00400693",
x"00d70463",
x"00478793",
x"00579713",
x"0037d793",
x"02075863",
x"00000793",
x"00100713",
x"f59ff06f",
x"00000793",
x"0ff00713",
x"f4dff06f",
x"004007b7",
x"0ff00713",
x"00000993",
x"f3dff06f",
x"00000793",
x"00000713",
x"f31ff06f",
x"008006b7",
x"fff68693",
x"ff010113",
x"00a6f633",
x"01755713",
x"00812423",
x"01f55413",
x"00361513",
x"0175d613",
x"00b6f6b3",
x"01212023",
x"00112623",
x"0ff77913",
x"00912223",
x"0ff67613",
x"0ff00713",
x"01f5d593",
x"00369793",
x"00e61463",
x"00079463",
x"0015c593",
x"40c906b3",
x"18859063",
x"08d05c63",
x"02061663",
x"02078063",
x"fff90693",
x"00069863",
x"00a787b3",
x"00100913",
x"04c0006f",
x"0ff00713",
x"00e91e63",
x"00050793",
x"10c0006f",
x"0ff00713",
x"fee90ae3",
x"04000737",
x"00e7e7b3",
x"01b00613",
x"00100713",
x"00d64e63",
x"02000613",
x"00d7d733",
x"40d606b3",
x"00d796b3",
x"00d036b3",
x"00d76733",
x"00a707b3",
x"00579713",
x"0c075663",
x"00190913",
x"0ff00713",
x"2ce90a63",
x"7e000737",
x"0017f693",
x"fff70713",
x"0017d793",
x"00e7f7b3",
x"00d7e7b3",
x"0a40006f",
x"06068663",
x"41260733",
x"02091063",
x"0c050863",
x"fff70693",
x"f60684e3",
x"0ff00593",
x"02b71063",
x"0ff00913",
x"07c0006f",
x"0ff00693",
x"fed60ae3",
x"040006b7",
x"00d56533",
x"00070693",
x"01b00593",
x"00100713",
x"00d5ce63",
x"02000713",
x"40d70733",
x"00e51733",
x"00d555b3",
x"00e03733",
x"00e5e733",
x"00e787b3",
x"00060913",
x"f69ff06f",
x"00190713",
x"0fe77693",
x"04069c63",
x"04091263",
x"02050263",
x"f00788e3",
x"00a787b3",
x"00579713",
x"00075a63",
x"fc000737",
x"fff70713",
x"00e7f7b3",
x"00100913",
x"0077f713",
x"20070a63",
x"00f7f713",
x"00400693",
x"20d70463",
x"00478793",
x"2000006f",
x"f60502e3",
x"16079663",
x"00050793",
x"f59ff06f",
x"0ff00693",
x"1ed70063",
x"00f507b3",
x"0017d793",
x"00070913",
x"fc1ff06f",
x"06d05e63",
x"06061263",
x"ea0782e3",
x"fff90693",
x"00069863",
x"40f507b3",
x"00100913",
x"0340006f",
x"0ff00713",
x"e8e904e3",
x"01b00613",
x"00100713",
x"00d64e63",
x"02000613",
x"00d7d733",
x"40d606b3",
x"00d796b3",
x"00d036b3",
x"00d76733",
x"40e507b3",
x"00579713",
x"f60754e3",
x"040004b7",
x"fff48493",
x"0097f4b3",
x"1080006f",
x"0ff00713",
x"e4e900e3",
x"04000737",
x"00e7e7b3",
x"fb1ff06f",
x"06068e63",
x"41260733",
x"02091663",
x"1a050e63",
x"fff70693",
x"00069863",
x"40a787b3",
x"00058413",
x"f7dff06f",
x"0ff00813",
x"03071063",
x"0ff00913",
x"19c0006f",
x"0ff00693",
x"fed60ae3",
x"040006b7",
x"00d56533",
x"00070693",
x"01b00813",
x"00100713",
x"00d84e63",
x"02000713",
x"40d70733",
x"00e51733",
x"00d55833",
x"00e03733",
x"00e86733",
x"40e787b3",
x"00060913",
x"00058413",
x"f5dff06f",
x"00190713",
x"0fe77713",
x"04071c63",
x"02091c63",
x"00051863",
x"12079e63",
x"00000413",
x"0c00006f",
x"d8078ae3",
x"40f50733",
x"00571693",
x"40a787b3",
x"1206c063",
x"00070793",
x"e80716e3",
x"00000793",
x"fd9ff06f",
x"ea0510e3",
x"00058413",
x"de079ce3",
x"00000413",
x"020007b7",
x"0ff00913",
x"0800006f",
x"40f504b3",
x"00549713",
x"04075463",
x"40a784b3",
x"00058413",
x"00048513",
x"338000ef",
x"ffb50513",
x"00a494b3",
x"03254e63",
x"41250533",
x"00150513",
x"02000713",
x"40a70733",
x"00a4d7b3",
x"00e494b3",
x"009034b3",
x"0097e7b3",
x"00000913",
x"e19ff06f",
x"fc0492e3",
x"00000793",
x"00000913",
x"f5dff06f",
x"fc0007b7",
x"fff78793",
x"40a90933",
x"00f4f7b3",
x"df5ff06f",
x"0ff00913",
x"00000793",
x"00579713",
x"00075e63",
x"00190913",
x"0ff00713",
x"06e90663",
x"fc000737",
x"fff70713",
x"00e7f7b3",
x"0ff00713",
x"0037d793",
x"00e91863",
x"00078663",
x"004007b7",
x"00000413",
x"00c12083",
x"01791713",
x"01f41513",
x"7f8006b7",
x"00812403",
x"00979793",
x"00d77733",
x"0097d793",
x"00f767b3",
x"00412483",
x"00012903",
x"00a7e533",
x"01010113",
x"00008067",
x"00070913",
x"00058413",
x"d71ff06f",
x"00000793",
x"fa1ff06f",
x"00800637",
x"01755713",
x"fff60793",
x"0ff77713",
x"07e00593",
x"00a7f7b3",
x"01f55693",
x"04e5d663",
x"09d00593",
x"00e5da63",
x"80000537",
x"fff50513",
x"00a68533",
x"00008067",
x"00c7e533",
x"09500793",
x"00e7dc63",
x"f6a70713",
x"00e51533",
x"02068063",
x"40a00533",
x"00008067",
x"09600793",
x"40e787b3",
x"00f55533",
x"fe9ff06f",
x"00000513",
x"00008067",
x"ff010113",
x"00112623",
x"00812423",
x"00912223",
x"00050793",
x"0e050063",
x"41f55713",
x"00a74433",
x"40e40433",
x"01f55493",
x"00040513",
x"1b4000ef",
x"09e00793",
x"40a787b3",
x"09600713",
x"04f74063",
x"00800713",
x"0ae50e63",
x"ff850513",
x"00a41433",
x"00941413",
x"00945413",
x"01779793",
x"00c12083",
x"0087e7b3",
x"00812403",
x"01f49513",
x"00a7e533",
x"00412483",
x"01010113",
x"00008067",
x"09900713",
x"06f75463",
x"00500713",
x"40a70733",
x"01b50693",
x"00e45733",
x"00d41433",
x"00803433",
x"00876733",
x"fc000437",
x"fff40413",
x"00777693",
x"00877433",
x"00068a63",
x"00f77713",
x"00400693",
x"00d70463",
x"00440413",
x"00541713",
x"00075c63",
x"fc0007b7",
x"fff78793",
x"00f47433",
x"09f00793",
x"40a787b3",
x"00345413",
x"f6dff06f",
x"ffb50713",
x"00e41733",
x"fb1ff06f",
x"00000493",
x"00000413",
x"f55ff06f",
x"09600793",
x"f4dff06f",
x"00050613",
x"00000513",
x"0015f693",
x"00068463",
x"00c50533",
x"0015d593",
x"00161613",
x"fe0596e3",
x"00008067",
x"06054063",
x"0605c663",
x"00058613",
x"00050593",
x"fff00513",
x"02060c63",
x"00100693",
x"00b67a63",
x"00c05863",
x"00161613",
x"00169693",
x"feb66ae3",
x"00000513",
x"00c5e663",
x"40c585b3",
x"00d56533",
x"0016d693",
x"00165613",
x"fe0696e3",
x"00008067",
x"00008293",
x"fb5ff0ef",
x"00058513",
x"00028067",
x"40a00533",
x"00b04863",
x"40b005b3",
x"f9dff06f",
x"40b005b3",
x"00008293",
x"f91ff0ef",
x"40a00533",
x"00028067",
x"00008293",
x"0005ca63",
x"00054c63",
x"f79ff0ef",
x"00058513",
x"00028067",
x"40b005b3",
x"fe0558e3",
x"40a00533",
x"f61ff0ef",
x"40b00533",
x"00028067",
x"000107b7",
x"02f57a63",
x"10053793",
x"0017b793",
x"00379793",
x"00002737",
x"02000693",
x"40f686b3",
x"00f55533",
x"20070793",
x"00a787b3",
x"0007c503",
x"40a68533",
x"00008067",
x"01000737",
x"01800793",
x"fce57ae3",
x"01000793",
x"fcdff06f",
x"000015c0",
x"00001648",
x"000015cc",
x"00001648",
x"000015d4",
x"00001648",
x"000015cc",
x"000015c0",
x"000015c0",
x"000015d4",
x"000015cc",
x"0000159c",
x"0000159c",
x"0000159c",
x"000015d4",
x"02020100",
x"03030303",
x"04040404",
x"04040404",
x"05050505",
x"05050505",
x"05050505",
x"05050505",
x"06060606",
x"06060606",
x"06060606",
x"06060606",
x"06060606",
x"06060606",
x"06060606",
x"06060606",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"07070707",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"08080808",
x"00000000",
x"80000184",
x"800001ec",
x"80000254",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000001",
x"00000000",
x"abcd330e",
x"e66d1234",
x"0005deec",
x"0000000b",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"7f800000",
x"42b17217",
x"c2cff1b5",
x"3fb8aa3b",
x"3f317180",
x"3717f7d1",
x"3331bb4c",
x"35ddea0e",
x"388ab355",
x"3b360b61",
x"3e2aaaab",
x"7149f2ca",
x"3f800000",
x"40000000",
x"0d800000",
x"10000000",
x"70000000",
x"bf800000",
x"3717f7d1",
x"b717f7d1",
x"3f317180",
x"bf317180",
x"3f000000",
x"bf000000",
x"80000000"
);

end neorv32_application_image;
